version https://git-lfs.github.com/spec/v1
oid sha256:b072267b8d5c6956711417e919e4e7b84fd66c4d786a800a227efd45a7cf838c
size 2141
