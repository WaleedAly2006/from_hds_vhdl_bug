version https://git-lfs.github.com/spec/v1
oid sha256:f105c05cdbde9230d59b79eb9eaa3d87cc3f43329f3f7c11f9f23389117230ff
size 13739
