version https://git-lfs.github.com/spec/v1
oid sha256:fc28d24084828b3dcb797fcf3269df027f11c2e216ed36073260e9c696a963c5
size 1480
