version https://git-lfs.github.com/spec/v1
oid sha256:364d1516908e5a4721e8fc569c7778ac1153a1343e244a2c6570b2d70f8fdc84
size 2849
