version https://git-lfs.github.com/spec/v1
oid sha256:91b53a2ee355500420f6b75b8597e67874931c367a582e466e78d2eb06de2006
size 9772
