version https://git-lfs.github.com/spec/v1
oid sha256:c07c928b48ec029057081eae6732774cbca1aa167b7f2efdf2fc3dae9ac06b39
size 2289
