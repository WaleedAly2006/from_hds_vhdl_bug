version https://git-lfs.github.com/spec/v1
oid sha256:0cf39d0b2a6f2f2a1ce0a4b9d13532b598a49994580066f0f6d4872d228c495a
size 6831
