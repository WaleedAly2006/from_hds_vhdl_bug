version https://git-lfs.github.com/spec/v1
oid sha256:cdc1e3098c97406f14a2157eec33ed5a43ecbd80fd50af58294df7c755bf925f
size 3534
