version https://git-lfs.github.com/spec/v1
oid sha256:72916290c917166eafa1fbdd73d05dad94d380e6d0c08809c351f6c7e98bb442
size 5959
